
module probes (
	source,
	probe);	

	output	[21:0]	source;
	input	[29:0]	probe;
endmodule
