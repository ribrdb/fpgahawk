// clocks.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module clocks (
		input  wire  clk_clk,             //           clk.clk
		output wire  pll_0_clk_100_clk,   // pll_0_clk_100.clk
		output wire  pll_0_clk_25_clk,    //  pll_0_clk_25.clk
		output wire  pll_0_clk_2_5_clk,   // pll_0_clk_2_5.clk
		output wire  pll_0_locked_export, //  pll_0_locked.export
		output wire  pll_1_locked_export, //  pll_1_locked.export
		output wire  pll_1_outclk0_clk,   // pll_1_outclk0.clk
		input  wire  reset_reset_n        //         reset.reset_n
	);

	clocks_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_clk_100_clk),   // outclk0.clk
		.outclk_1 (pll_0_clk_25_clk),    // outclk1.clk
		.outclk_2 (pll_0_clk_2_5_clk),   // outclk2.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	clocks_pll_1 pll_1 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_1_outclk0_clk),   // outclk0.clk
		.locked   (pll_1_locked_export)  //  locked.export
	);

endmodule
